module dp_tb;

    initial begin

    end

endmodule