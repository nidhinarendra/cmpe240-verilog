module dp();

    reg [7:0] memA [7:0];
    reg [7:0] memb [7:0];

endmodule