module mem_transfer();

endmodule