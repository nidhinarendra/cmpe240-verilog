module counter();

endmodule

module dreg();

endmodule

module comparator();

endmodule

module adder();

endmodule

module sub();

endmodule

module mux2to1();

endmodule