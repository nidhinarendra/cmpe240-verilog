module cu_tb;

initial begin


end

endmodule