module mem_transfer_tb;

    initial begin
    
    end
endmodule